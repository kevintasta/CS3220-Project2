library verilog;
use verilog.vl_types.all;
entity TestSignExtension is
end TestSignExtension;
