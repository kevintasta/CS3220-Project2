library verilog;
use verilog.vl_types.all;
entity TestBranchPicker is
end TestBranchPicker;
