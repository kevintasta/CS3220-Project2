library verilog;
use verilog.vl_types.all;
entity TestProject2 is
end TestProject2;
