library verilog;
use verilog.vl_types.all;
entity TestAdder is
end TestAdder;
