library verilog;
use verilog.vl_types.all;
entity TestMultiplexer is
end TestMultiplexer;
