library verilog;
use verilog.vl_types.all;
entity TestRegister is
end TestRegister;
