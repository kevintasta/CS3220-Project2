library verilog;
use verilog.vl_types.all;
entity TestLeftShift is
end TestLeftShift;
